library IEEE;
use IEEE.std_logic_1164.all;
----------------------------------------------
ENTITY ss_counter IS
	PORT (clk, toggle: IN std_logic;
			count: OUT INTEGER RANGE 0 TO 9);
END ENTITY;
----------------------------------------------
ARCHITECTURE ss_counter OF ss_counter IS
SIGNAL temp: INTEGER RANGE 0 TO 10;
BEGIN
	PROCESS(clk, toggle)
	BEGIN
		IF (toggle = '0') THEN
			IF (clk'EVENt AND clk='1') THEN
				IF (temp = 9) THEN
					temp <= 0;
				ELSE
					temp <= temp + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	count <= temp;
END ARCHITECTURE;
----------------------------------------------
